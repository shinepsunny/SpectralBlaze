
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "df_loop_interface.svh"
`include "df_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_fwd_fft.c_ifmap_patch_st_U.if_read;
    assign fifo_intf_1.wr_en = AESL_inst_fwd_fft.c_ifmap_patch_st_U.if_write;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.c_ifmap_patch_st_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.c_ifmap_patch_st_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_fwd_fft.ctrl1_reg_c21_U.if_read;
    assign fifo_intf_2.wr_en = AESL_inst_fwd_fft.ctrl1_reg_c21_U.if_write;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl1_reg_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ctrl1_reg_c21_blk_n);
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_fwd_fft.ctrl2_reg_c26_U.if_read;
    assign fifo_intf_3.wr_en = AESL_inst_fwd_fft.ctrl2_reg_c26_U.if_write;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl2_reg_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ctrl2_reg_c26_blk_n);
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_fwd_fft.layer1_reg_c31_U.if_read;
    assign fifo_intf_4.wr_en = AESL_inst_fwd_fft.layer1_reg_c31_U.if_write;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.layer1_reg_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_fwd_fft.Mem_Patch_Gen_U0.layer1_reg_c31_blk_n);
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_fwd_fft.c_ifmap_col_op_st_U.if_read;
    assign fifo_intf_5.wr_en = AESL_inst_fwd_fft.c_ifmap_col_op_st_U.if_write;
    assign fifo_intf_5.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.c_row_op_trans_st_blk_n);
    assign fifo_intf_5.fifo_wr_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.c_ifmap_col_op_st_blk_n);
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_fwd_fft.ctrl1_reg_c20_U.if_read;
    assign fifo_intf_6.wr_en = AESL_inst_fwd_fft.ctrl1_reg_c20_U.if_write;
    assign fifo_intf_6.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_R_U0.ctrl1_reg_blk_n);
    assign fifo_intf_6.fifo_wr_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl1_reg_c20_blk_n);
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_fwd_fft.ctrl2_reg_c25_U.if_read;
    assign fifo_intf_7.wr_en = AESL_inst_fwd_fft.ctrl2_reg_c25_U.if_write;
    assign fifo_intf_7.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_R_U0.ctrl2_reg_blk_n);
    assign fifo_intf_7.fifo_wr_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl2_reg_c25_blk_n);
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_fwd_fft.layer1_reg_c30_U.if_read;
    assign fifo_intf_8.wr_en = AESL_inst_fwd_fft.layer1_reg_c30_U.if_write;
    assign fifo_intf_8.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_R_U0.layer1_reg_blk_n);
    assign fifo_intf_8.fifo_wr_block = ~(AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.layer1_reg_c30_blk_n);
    assign fifo_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_fwd_fft.c_fft_row_op_st_U.if_read;
    assign fifo_intf_9.wr_en = AESL_inst_fwd_fft.c_fft_row_op_st_U.if_write;
    assign fifo_intf_9.fifo_rd_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.c_fft_row_op_st_blk_n);
    assign fifo_intf_9.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.c_fft_col_op_st_blk_n);
    assign fifo_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_fwd_fft.ctrl1_reg_c19_U.if_read;
    assign fifo_intf_10.wr_en = AESL_inst_fwd_fft.ctrl1_reg_c19_U.if_write;
    assign fifo_intf_10.fifo_rd_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl1_reg_blk_n);
    assign fifo_intf_10.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_R_U0.ctrl1_reg_c19_blk_n);
    assign fifo_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_fwd_fft.ctrl2_reg_c24_U.if_read;
    assign fifo_intf_11.wr_en = AESL_inst_fwd_fft.ctrl2_reg_c24_U.if_write;
    assign fifo_intf_11.fifo_rd_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl2_reg_blk_n);
    assign fifo_intf_11.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_R_U0.ctrl2_reg_c24_blk_n);
    assign fifo_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_fwd_fft.layer1_reg_c29_U.if_read;
    assign fifo_intf_12.wr_en = AESL_inst_fwd_fft.layer1_reg_c29_U.if_write;
    assign fifo_intf_12.fifo_rd_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.layer1_reg_blk_n);
    assign fifo_intf_12.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_R_U0.layer1_reg_c29_blk_n);
    assign fifo_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c6_channel_U.if_read;
    assign fifo_intf_13.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c6_channel_U.if_write;
    assign fifo_intf_13.fifo_rd_block = 0;
    assign fifo_intf_13.fifo_wr_block = 0;
    assign fifo_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c5_channel_U.if_read;
    assign fifo_intf_14.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c5_channel_U.if_write;
    assign fifo_intf_14.fifo_rd_block = 0;
    assign fifo_intf_14.fifo_wr_block = 0;
    assign fifo_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c4_channel_U.if_read;
    assign fifo_intf_15.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c4_channel_U.if_write;
    assign fifo_intf_15.fifo_rd_block = 0;
    assign fifo_intf_15.fifo_wr_block = 0;
    assign fifo_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c3_channel_U.if_read;
    assign fifo_intf_16.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c3_channel_U.if_write;
    assign fifo_intf_16.fifo_rd_block = 0;
    assign fifo_intf_16.fifo_wr_block = 0;
    assign fifo_intf_16.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c2_channel_U.if_read;
    assign fifo_intf_17.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c2_channel_U.if_write;
    assign fifo_intf_17.fifo_rd_block = 0;
    assign fifo_intf_17.fifo_wr_block = 0;
    assign fifo_intf_17.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c1_channel_U.if_read;
    assign fifo_intf_18.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c1_channel_U.if_write;
    assign fifo_intf_18.fifo_rd_block = 0;
    assign fifo_intf_18.fifo_wr_block = 0;
    assign fifo_intf_18.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c_channel_U.if_read;
    assign fifo_intf_19.wr_en = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ctrl1_reg_c_channel_U.if_write;
    assign fifo_intf_19.fifo_rd_block = 0;
    assign fifo_intf_19.fifo_wr_block = 0;
    assign fifo_intf_19.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_fwd_fft.c_row_op_st_U.if_read;
    assign fifo_intf_20.wr_en = AESL_inst_fwd_fft.c_row_op_st_U.if_write;
    assign fifo_intf_20.fifo_rd_block = ~(AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.c_row_op_st_blk_n);
    assign fifo_intf_20.fifo_wr_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.c_row_op_st_blk_n & AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.c_row_op_st_blk_n);
    assign fifo_intf_20.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_fwd_fft.ctrl1_reg_c18_U.if_read;
    assign fifo_intf_21.wr_en = AESL_inst_fwd_fft.ctrl1_reg_c18_U.if_write;
    assign fifo_intf_21.fifo_rd_block = ~(AESL_inst_fwd_fft.Transpose_U0.ctrl1_reg_blk_n);
    assign fifo_intf_21.fifo_wr_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl1_reg_c18_blk_n);
    assign fifo_intf_21.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_fwd_fft.ctrl2_reg_c23_U.if_read;
    assign fifo_intf_22.wr_en = AESL_inst_fwd_fft.ctrl2_reg_c23_U.if_write;
    assign fifo_intf_22.fifo_rd_block = ~(AESL_inst_fwd_fft.Transpose_U0.ctrl2_reg_blk_n);
    assign fifo_intf_22.fifo_wr_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl2_reg_c23_blk_n);
    assign fifo_intf_22.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_fwd_fft.layer1_reg_c28_U.if_read;
    assign fifo_intf_23.wr_en = AESL_inst_fwd_fft.layer1_reg_c28_U.if_write;
    assign fifo_intf_23.fifo_rd_block = ~(AESL_inst_fwd_fft.Transpose_U0.layer1_reg_blk_n);
    assign fifo_intf_23.fifo_wr_block = ~(AESL_inst_fwd_fft.Row_Wise_Synch_U0.layer1_reg_c28_blk_n);
    assign fifo_intf_23.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_fwd_fft.c_row_op_trans_st_U.if_read;
    assign fifo_intf_24.wr_en = AESL_inst_fwd_fft.c_row_op_trans_st_U.if_write;
    assign fifo_intf_24.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.c_row_op_trans_st_blk_n);
    assign fifo_intf_24.fifo_wr_block = ~(AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.c_row_op_trans_st_blk_n);
    assign fifo_intf_24.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_fwd_fft.ctrl1_reg_c17_U.if_read;
    assign fifo_intf_25.wr_en = AESL_inst_fwd_fft.ctrl1_reg_c17_U.if_write;
    assign fifo_intf_25.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_C_U0.ctrl1_reg_blk_n);
    assign fifo_intf_25.fifo_wr_block = ~(AESL_inst_fwd_fft.Transpose_U0.ctrl1_reg_c17_blk_n);
    assign fifo_intf_25.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_fwd_fft.ctrl2_reg_c22_U.if_read;
    assign fifo_intf_26.wr_en = AESL_inst_fwd_fft.ctrl2_reg_c22_U.if_write;
    assign fifo_intf_26.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_C_U0.ctrl2_reg_blk_n);
    assign fifo_intf_26.fifo_wr_block = ~(AESL_inst_fwd_fft.Transpose_U0.ctrl2_reg_c22_blk_n);
    assign fifo_intf_26.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_fwd_fft.layer1_reg_c27_U.if_read;
    assign fifo_intf_27.wr_en = AESL_inst_fwd_fft.layer1_reg_c27_U.if_write;
    assign fifo_intf_27.fifo_rd_block = ~(AESL_inst_fwd_fft.FFT_C_U0.layer1_reg_blk_n);
    assign fifo_intf_27.fifo_wr_block = ~(AESL_inst_fwd_fft.Transpose_U0.layer1_reg_c27_blk_n);
    assign fifo_intf_27.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ctrl1_reg_c_channel1_U.if_read;
    assign fifo_intf_28.wr_en = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ctrl1_reg_c_channel1_U.if_write;
    assign fifo_intf_28.fifo_rd_block = 0;
    assign fifo_intf_28.fifo_wr_block = 0;
    assign fifo_intf_28.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_fwd_fft.c_fft_col_op_st_U.if_read;
    assign fifo_intf_29.wr_en = AESL_inst_fwd_fft.c_fft_col_op_st_U.if_write;
    assign fifo_intf_29.fifo_rd_block = ~(AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.c_fft_col_op_st_blk_n);
    assign fifo_intf_29.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.c_fft_col_op_st_blk_n);
    assign fifo_intf_29.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_fwd_fft.ctrl1_reg_c_U.if_read;
    assign fifo_intf_30.wr_en = AESL_inst_fwd_fft.ctrl1_reg_c_U.if_write;
    assign fifo_intf_30.fifo_rd_block = ~(AESL_inst_fwd_fft.Mem_patch_Wr_U0.ctrl1_reg_blk_n);
    assign fifo_intf_30.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_C_U0.ctrl1_reg_c_blk_n);
    assign fifo_intf_30.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_fwd_fft.ctrl2_reg_c_U.if_read;
    assign fifo_intf_31.wr_en = AESL_inst_fwd_fft.ctrl2_reg_c_U.if_write;
    assign fifo_intf_31.fifo_rd_block = ~(AESL_inst_fwd_fft.Mem_patch_Wr_U0.ctrl2_reg_blk_n);
    assign fifo_intf_31.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_C_U0.ctrl2_reg_c_blk_n);
    assign fifo_intf_31.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_fwd_fft.layer1_reg_c_U.if_read;
    assign fifo_intf_32.wr_en = AESL_inst_fwd_fft.layer1_reg_c_U.if_write;
    assign fifo_intf_32.fifo_rd_block = ~(AESL_inst_fwd_fft.Mem_patch_Wr_U0.layer1_reg_blk_n);
    assign fifo_intf_32.fifo_wr_block = ~(AESL_inst_fwd_fft.FFT_C_U0.layer1_reg_c_blk_n);
    assign fifo_intf_32.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c6_channel_U.if_read;
    assign fifo_intf_33.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c6_channel_U.if_write;
    assign fifo_intf_33.fifo_rd_block = 0;
    assign fifo_intf_33.fifo_wr_block = 0;
    assign fifo_intf_33.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c5_channel_U.if_read;
    assign fifo_intf_34.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c5_channel_U.if_write;
    assign fifo_intf_34.fifo_rd_block = 0;
    assign fifo_intf_34.fifo_wr_block = 0;
    assign fifo_intf_34.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;
    df_fifo_intf fifo_intf_35(clock,reset);
    assign fifo_intf_35.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c4_channel_U.if_read;
    assign fifo_intf_35.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c4_channel_U.if_write;
    assign fifo_intf_35.fifo_rd_block = 0;
    assign fifo_intf_35.fifo_wr_block = 0;
    assign fifo_intf_35.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_35;
    csv_file_dump cstatus_csv_dumper_35;
    df_fifo_monitor fifo_monitor_35;
    df_fifo_intf fifo_intf_36(clock,reset);
    assign fifo_intf_36.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c3_channel_U.if_read;
    assign fifo_intf_36.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c3_channel_U.if_write;
    assign fifo_intf_36.fifo_rd_block = 0;
    assign fifo_intf_36.fifo_wr_block = 0;
    assign fifo_intf_36.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_36;
    csv_file_dump cstatus_csv_dumper_36;
    df_fifo_monitor fifo_monitor_36;
    df_fifo_intf fifo_intf_37(clock,reset);
    assign fifo_intf_37.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c2_channel_U.if_read;
    assign fifo_intf_37.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c2_channel_U.if_write;
    assign fifo_intf_37.fifo_rd_block = 0;
    assign fifo_intf_37.fifo_wr_block = 0;
    assign fifo_intf_37.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_37;
    csv_file_dump cstatus_csv_dumper_37;
    df_fifo_monitor fifo_monitor_37;
    df_fifo_intf fifo_intf_38(clock,reset);
    assign fifo_intf_38.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c1_channel_U.if_read;
    assign fifo_intf_38.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c1_channel_U.if_write;
    assign fifo_intf_38.fifo_rd_block = 0;
    assign fifo_intf_38.fifo_wr_block = 0;
    assign fifo_intf_38.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_38;
    csv_file_dump cstatus_csv_dumper_38;
    df_fifo_monitor fifo_monitor_38;
    df_fifo_intf fifo_intf_39(clock,reset);
    assign fifo_intf_39.rd_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c_channel_U.if_read;
    assign fifo_intf_39.wr_en = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ctrl1_reg_c_channel_U.if_write;
    assign fifo_intf_39.fifo_rd_block = 0;
    assign fifo_intf_39.fifo_wr_block = 0;
    assign fifo_intf_39.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_39;
    csv_file_dump cstatus_csv_dumper_39;
    df_fifo_monitor fifo_monitor_39;
    df_fifo_intf fifo_intf_40(clock,reset);
    assign fifo_intf_40.rd_en = AESL_inst_fwd_fft.out_c_channel_U.if_read;
    assign fifo_intf_40.wr_en = AESL_inst_fwd_fft.out_c_channel_U.if_write;
    assign fifo_intf_40.fifo_rd_block = 0;
    assign fifo_intf_40.fifo_wr_block = 0;
    assign fifo_intf_40.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_40;
    csv_file_dump cstatus_csv_dumper_40;
    df_fifo_monitor fifo_monitor_40;
    df_fifo_intf fifo_intf_41(clock,reset);
    assign fifo_intf_41.rd_en = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.fft_out_c_channel_U.if_read;
    assign fifo_intf_41.wr_en = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.fft_out_c_channel_U.if_write;
    assign fifo_intf_41.fifo_rd_block = 0;
    assign fifo_intf_41.fifo_wr_block = 0;
    assign fifo_intf_41.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_41;
    csv_file_dump cstatus_csv_dumper_41;
    df_fifo_monitor fifo_monitor_41;
    df_fifo_intf fifo_intf_42(clock,reset);
    assign fifo_intf_42.rd_en = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ctrl1_reg_c_channel1_U.if_read;
    assign fifo_intf_42.wr_en = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ctrl1_reg_c_channel1_U.if_write;
    assign fifo_intf_42.fifo_rd_block = 0;
    assign fifo_intf_42.fifo_wr_block = 0;
    assign fifo_intf_42.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_42;
    csv_file_dump cstatus_csv_dumper_42;
    df_fifo_monitor fifo_monitor_42;

    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_fwd_fft.entry_proc47_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_fwd_fft.entry_proc47_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_fwd_fft.entry_proc47_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_fwd_fft.entry_proc47_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_fwd_fft.entry_proc47_U0.ap_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.real_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0 | ~AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.c_ifmap_patch_st_blk_n | ~AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ctrl1_reg_c21_blk_n | ~AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ctrl2_reg_c26_blk_n | ~AESL_inst_fwd_fft.Mem_Patch_Gen_U0.layer1_reg_c31_blk_n;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.real_start;
    assign process_intf_3.pin_stall = 1'b0 | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.c_ifmap_patch_st_blk_n | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl1_reg_blk_n | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl2_reg_blk_n | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.layer1_reg_blk_n;
    assign process_intf_3.pout_stall = 1'b0 | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.c_ifmap_col_op_st_blk_n | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl1_reg_c20_blk_n | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.ctrl2_reg_c25_blk_n | ~AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.layer1_reg_c30_blk_n;
    assign process_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_fwd_fft.FFT_R_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_fwd_fft.FFT_R_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_fwd_fft.FFT_R_U0.real_start;
    assign process_intf_4.pin_stall = 1'b0 | ~AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.c_row_op_trans_st_blk_n | ~AESL_inst_fwd_fft.FFT_R_U0.ctrl1_reg_blk_n | ~AESL_inst_fwd_fft.FFT_R_U0.ctrl2_reg_blk_n | ~AESL_inst_fwd_fft.FFT_R_U0.layer1_reg_blk_n;
    assign process_intf_4.pout_stall = 1'b0 | ~AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.c_fft_col_op_st_blk_n | ~AESL_inst_fwd_fft.FFT_R_U0.ctrl1_reg_c19_blk_n | ~AESL_inst_fwd_fft.FFT_R_U0.ctrl2_reg_c24_blk_n | ~AESL_inst_fwd_fft.FFT_R_U0.layer1_reg_c29_blk_n;
    assign process_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_start;
    assign process_intf_5.pin_stall = 1'b0;
    assign process_intf_5.pout_stall = 1'b0;
    assign process_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;
    df_process_intf process_intf_6(clock,reset);
    assign process_intf_6.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_start;
    assign process_intf_6.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_ready;
    assign process_intf_6.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_done;
    assign process_intf_6.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_continue;
    assign process_intf_6.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_start;
    assign process_intf_6.pin_stall = 1'b0;
    assign process_intf_6.pout_stall = 1'b0;
    assign process_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_6;
    csv_file_dump pstatus_csv_dumper_6;
    df_process_monitor process_monitor_6;
    df_process_intf process_intf_7(clock,reset);
    assign process_intf_7.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.ap_start;
    assign process_intf_7.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.ap_ready;
    assign process_intf_7.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.ap_done;
    assign process_intf_7.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.ap_continue;
    assign process_intf_7.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.ap_start;
    assign process_intf_7.pin_stall = 1'b0;
    assign process_intf_7.pout_stall = 1'b0;
    assign process_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_7;
    csv_file_dump pstatus_csv_dumper_7;
    df_process_monitor process_monitor_7;
    df_process_intf process_intf_8(clock,reset);
    assign process_intf_8.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.ap_start;
    assign process_intf_8.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.ap_ready;
    assign process_intf_8.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.ap_done;
    assign process_intf_8.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.ap_continue;
    assign process_intf_8.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.ap_start;
    assign process_intf_8.pin_stall = 1'b0;
    assign process_intf_8.pout_stall = 1'b0;
    assign process_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_8;
    csv_file_dump pstatus_csv_dumper_8;
    df_process_monitor process_monitor_8;
    df_process_intf process_intf_9(clock,reset);
    assign process_intf_9.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.ap_start;
    assign process_intf_9.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.ap_ready;
    assign process_intf_9.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.ap_done;
    assign process_intf_9.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.ap_continue;
    assign process_intf_9.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.ap_start;
    assign process_intf_9.pin_stall = 1'b0;
    assign process_intf_9.pout_stall = 1'b0;
    assign process_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_9;
    csv_file_dump pstatus_csv_dumper_9;
    df_process_monitor process_monitor_9;
    df_process_intf process_intf_10(clock,reset);
    assign process_intf_10.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.ap_start;
    assign process_intf_10.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.ap_ready;
    assign process_intf_10.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.ap_done;
    assign process_intf_10.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.ap_continue;
    assign process_intf_10.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.ap_start;
    assign process_intf_10.pin_stall = 1'b0;
    assign process_intf_10.pout_stall = 1'b0;
    assign process_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_10;
    csv_file_dump pstatus_csv_dumper_10;
    df_process_monitor process_monitor_10;
    df_process_intf process_intf_11(clock,reset);
    assign process_intf_11.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.ap_start;
    assign process_intf_11.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.ap_ready;
    assign process_intf_11.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.ap_done;
    assign process_intf_11.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.ap_continue;
    assign process_intf_11.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.ap_start;
    assign process_intf_11.pin_stall = 1'b0;
    assign process_intf_11.pout_stall = 1'b0;
    assign process_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_11;
    csv_file_dump pstatus_csv_dumper_11;
    df_process_monitor process_monitor_11;
    df_process_intf process_intf_12(clock,reset);
    assign process_intf_12.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.ap_start;
    assign process_intf_12.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.ap_ready;
    assign process_intf_12.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.ap_done;
    assign process_intf_12.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.ap_continue;
    assign process_intf_12.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.ap_start;
    assign process_intf_12.pin_stall = 1'b0;
    assign process_intf_12.pout_stall = 1'b0;
    assign process_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_12;
    csv_file_dump pstatus_csv_dumper_12;
    df_process_monitor process_monitor_12;
    df_process_intf process_intf_13(clock,reset);
    assign process_intf_13.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_start;
    assign process_intf_13.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_ready;
    assign process_intf_13.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_done;
    assign process_intf_13.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_continue;
    assign process_intf_13.real_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_start;
    assign process_intf_13.pin_stall = 1'b0;
    assign process_intf_13.pout_stall = 1'b0;
    assign process_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_13;
    csv_file_dump pstatus_csv_dumper_13;
    df_process_monitor process_monitor_13;
    df_process_intf process_intf_14(clock,reset);
    assign process_intf_14.ap_start = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_start;
    assign process_intf_14.ap_ready = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_ready;
    assign process_intf_14.ap_done = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_done;
    assign process_intf_14.ap_continue = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_continue;
    assign process_intf_14.real_start = AESL_inst_fwd_fft.Row_Wise_Synch_U0.real_start;
    assign process_intf_14.pin_stall = 1'b0 | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.c_fft_row_op_st_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl1_reg_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl2_reg_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.layer1_reg_blk_n;
    assign process_intf_14.pout_stall = 1'b0 | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.c_row_op_st_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.c_row_op_st_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl1_reg_c18_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.ctrl2_reg_c23_blk_n | ~AESL_inst_fwd_fft.Row_Wise_Synch_U0.layer1_reg_c28_blk_n;
    assign process_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_14;
    csv_file_dump pstatus_csv_dumper_14;
    df_process_monitor process_monitor_14;
    df_process_intf process_intf_15(clock,reset);
    assign process_intf_15.ap_start = AESL_inst_fwd_fft.Transpose_U0.ap_start;
    assign process_intf_15.ap_ready = AESL_inst_fwd_fft.Transpose_U0.ap_ready;
    assign process_intf_15.ap_done = AESL_inst_fwd_fft.Transpose_U0.ap_done;
    assign process_intf_15.ap_continue = AESL_inst_fwd_fft.Transpose_U0.ap_continue;
    assign process_intf_15.real_start = AESL_inst_fwd_fft.Transpose_U0.real_start;
    assign process_intf_15.pin_stall = 1'b0 | ~AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.c_row_op_st_blk_n | ~AESL_inst_fwd_fft.Transpose_U0.ctrl1_reg_blk_n | ~AESL_inst_fwd_fft.Transpose_U0.ctrl2_reg_blk_n | ~AESL_inst_fwd_fft.Transpose_U0.layer1_reg_blk_n;
    assign process_intf_15.pout_stall = 1'b0 | ~AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.c_row_op_trans_st_blk_n | ~AESL_inst_fwd_fft.Transpose_U0.ctrl1_reg_c17_blk_n | ~AESL_inst_fwd_fft.Transpose_U0.ctrl2_reg_c22_blk_n | ~AESL_inst_fwd_fft.Transpose_U0.layer1_reg_c27_blk_n;
    assign process_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_15;
    csv_file_dump pstatus_csv_dumper_15;
    df_process_monitor process_monitor_15;
    df_process_intf process_intf_16(clock,reset);
    assign process_intf_16.ap_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_start;
    assign process_intf_16.ap_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_ready;
    assign process_intf_16.ap_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_done;
    assign process_intf_16.ap_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_continue;
    assign process_intf_16.real_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_start;
    assign process_intf_16.pin_stall = 1'b0;
    assign process_intf_16.pout_stall = 1'b0;
    assign process_intf_16.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_16;
    csv_file_dump pstatus_csv_dumper_16;
    df_process_monitor process_monitor_16;
    df_process_intf process_intf_17(clock,reset);
    assign process_intf_17.ap_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_start;
    assign process_intf_17.ap_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_ready;
    assign process_intf_17.ap_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_done;
    assign process_intf_17.ap_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_continue;
    assign process_intf_17.real_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_start;
    assign process_intf_17.pin_stall = 1'b0;
    assign process_intf_17.pout_stall = 1'b0;
    assign process_intf_17.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_17;
    csv_file_dump pstatus_csv_dumper_17;
    df_process_monitor process_monitor_17;
    df_process_intf process_intf_18(clock,reset);
    assign process_intf_18.ap_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_start;
    assign process_intf_18.ap_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_ready;
    assign process_intf_18.ap_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_done;
    assign process_intf_18.ap_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_continue;
    assign process_intf_18.real_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_start;
    assign process_intf_18.pin_stall = 1'b0;
    assign process_intf_18.pout_stall = 1'b0;
    assign process_intf_18.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_18;
    csv_file_dump pstatus_csv_dumper_18;
    df_process_monitor process_monitor_18;
    df_process_intf process_intf_19(clock,reset);
    assign process_intf_19.ap_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_start;
    assign process_intf_19.ap_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_ready;
    assign process_intf_19.ap_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_done;
    assign process_intf_19.ap_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_continue;
    assign process_intf_19.real_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_start;
    assign process_intf_19.pin_stall = 1'b0;
    assign process_intf_19.pout_stall = 1'b0;
    assign process_intf_19.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_19;
    csv_file_dump pstatus_csv_dumper_19;
    df_process_monitor process_monitor_19;
    df_process_intf process_intf_20(clock,reset);
    assign process_intf_20.ap_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_start;
    assign process_intf_20.ap_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_ready;
    assign process_intf_20.ap_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_done;
    assign process_intf_20.ap_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_continue;
    assign process_intf_20.real_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_start;
    assign process_intf_20.pin_stall = 1'b0;
    assign process_intf_20.pout_stall = 1'b0;
    assign process_intf_20.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_20;
    csv_file_dump pstatus_csv_dumper_20;
    df_process_monitor process_monitor_20;
    df_process_intf process_intf_21(clock,reset);
    assign process_intf_21.ap_start = AESL_inst_fwd_fft.FFT_C_U0.ap_start;
    assign process_intf_21.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.ap_ready;
    assign process_intf_21.ap_done = AESL_inst_fwd_fft.FFT_C_U0.ap_done;
    assign process_intf_21.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.ap_continue;
    assign process_intf_21.real_start = AESL_inst_fwd_fft.FFT_C_U0.ap_start;
    assign process_intf_21.pin_stall = 1'b0 | ~AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.c_row_op_trans_st_blk_n | ~AESL_inst_fwd_fft.FFT_C_U0.ctrl1_reg_blk_n | ~AESL_inst_fwd_fft.FFT_C_U0.ctrl2_reg_blk_n | ~AESL_inst_fwd_fft.FFT_C_U0.layer1_reg_blk_n;
    assign process_intf_21.pout_stall = 1'b0 | ~AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.c_fft_col_op_st_blk_n | ~AESL_inst_fwd_fft.FFT_C_U0.ctrl1_reg_c_blk_n | ~AESL_inst_fwd_fft.FFT_C_U0.ctrl2_reg_c_blk_n | ~AESL_inst_fwd_fft.FFT_C_U0.layer1_reg_c_blk_n;
    assign process_intf_21.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_21;
    csv_file_dump pstatus_csv_dumper_21;
    df_process_monitor process_monitor_21;
    df_process_intf process_intf_22(clock,reset);
    assign process_intf_22.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_start;
    assign process_intf_22.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_ready;
    assign process_intf_22.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_done;
    assign process_intf_22.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_continue;
    assign process_intf_22.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_start;
    assign process_intf_22.pin_stall = 1'b0;
    assign process_intf_22.pout_stall = 1'b0;
    assign process_intf_22.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_22;
    csv_file_dump pstatus_csv_dumper_22;
    df_process_monitor process_monitor_22;
    df_process_intf process_intf_23(clock,reset);
    assign process_intf_23.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_start;
    assign process_intf_23.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_ready;
    assign process_intf_23.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_done;
    assign process_intf_23.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_continue;
    assign process_intf_23.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_start;
    assign process_intf_23.pin_stall = 1'b0;
    assign process_intf_23.pout_stall = 1'b0;
    assign process_intf_23.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_23;
    csv_file_dump pstatus_csv_dumper_23;
    df_process_monitor process_monitor_23;
    df_process_intf process_intf_24(clock,reset);
    assign process_intf_24.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.ap_start;
    assign process_intf_24.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.ap_ready;
    assign process_intf_24.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.ap_done;
    assign process_intf_24.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.ap_continue;
    assign process_intf_24.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.ap_start;
    assign process_intf_24.pin_stall = 1'b0;
    assign process_intf_24.pout_stall = 1'b0;
    assign process_intf_24.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_24;
    csv_file_dump pstatus_csv_dumper_24;
    df_process_monitor process_monitor_24;
    df_process_intf process_intf_25(clock,reset);
    assign process_intf_25.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.ap_start;
    assign process_intf_25.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.ap_ready;
    assign process_intf_25.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.ap_done;
    assign process_intf_25.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.ap_continue;
    assign process_intf_25.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.ap_start;
    assign process_intf_25.pin_stall = 1'b0;
    assign process_intf_25.pout_stall = 1'b0;
    assign process_intf_25.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_25;
    csv_file_dump pstatus_csv_dumper_25;
    df_process_monitor process_monitor_25;
    df_process_intf process_intf_26(clock,reset);
    assign process_intf_26.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.ap_start;
    assign process_intf_26.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.ap_ready;
    assign process_intf_26.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.ap_done;
    assign process_intf_26.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.ap_continue;
    assign process_intf_26.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.ap_start;
    assign process_intf_26.pin_stall = 1'b0;
    assign process_intf_26.pout_stall = 1'b0;
    assign process_intf_26.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_26;
    csv_file_dump pstatus_csv_dumper_26;
    df_process_monitor process_monitor_26;
    df_process_intf process_intf_27(clock,reset);
    assign process_intf_27.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.ap_start;
    assign process_intf_27.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.ap_ready;
    assign process_intf_27.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.ap_done;
    assign process_intf_27.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.ap_continue;
    assign process_intf_27.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.ap_start;
    assign process_intf_27.pin_stall = 1'b0;
    assign process_intf_27.pout_stall = 1'b0;
    assign process_intf_27.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_27;
    csv_file_dump pstatus_csv_dumper_27;
    df_process_monitor process_monitor_27;
    df_process_intf process_intf_28(clock,reset);
    assign process_intf_28.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.ap_start;
    assign process_intf_28.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.ap_ready;
    assign process_intf_28.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.ap_done;
    assign process_intf_28.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.ap_continue;
    assign process_intf_28.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.ap_start;
    assign process_intf_28.pin_stall = 1'b0;
    assign process_intf_28.pout_stall = 1'b0;
    assign process_intf_28.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_28;
    csv_file_dump pstatus_csv_dumper_28;
    df_process_monitor process_monitor_28;
    df_process_intf process_intf_29(clock,reset);
    assign process_intf_29.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.ap_start;
    assign process_intf_29.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.ap_ready;
    assign process_intf_29.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.ap_done;
    assign process_intf_29.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.ap_continue;
    assign process_intf_29.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.ap_start;
    assign process_intf_29.pin_stall = 1'b0;
    assign process_intf_29.pout_stall = 1'b0;
    assign process_intf_29.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_29;
    csv_file_dump pstatus_csv_dumper_29;
    df_process_monitor process_monitor_29;
    df_process_intf process_intf_30(clock,reset);
    assign process_intf_30.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_start;
    assign process_intf_30.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_ready;
    assign process_intf_30.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_done;
    assign process_intf_30.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_continue;
    assign process_intf_30.real_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_start;
    assign process_intf_30.pin_stall = 1'b0;
    assign process_intf_30.pout_stall = 1'b0;
    assign process_intf_30.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_30;
    csv_file_dump pstatus_csv_dumper_30;
    df_process_monitor process_monitor_30;
    df_process_intf process_intf_31(clock,reset);
    assign process_intf_31.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.ap_start;
    assign process_intf_31.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.ap_ready;
    assign process_intf_31.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.ap_done;
    assign process_intf_31.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.ap_continue;
    assign process_intf_31.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.ap_start;
    assign process_intf_31.pin_stall = 1'b0 | ~AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.c_fft_col_op_st_blk_n | ~AESL_inst_fwd_fft.Mem_patch_Wr_U0.ctrl1_reg_blk_n | ~AESL_inst_fwd_fft.Mem_patch_Wr_U0.ctrl2_reg_blk_n | ~AESL_inst_fwd_fft.Mem_patch_Wr_U0.layer1_reg_blk_n;
    assign process_intf_31.pout_stall = 1'b0;
    assign process_intf_31.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_31;
    csv_file_dump pstatus_csv_dumper_31;
    df_process_monitor process_monitor_31;
    df_process_intf process_intf_32(clock,reset);
    assign process_intf_32.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_start;
    assign process_intf_32.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_ready;
    assign process_intf_32.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_done;
    assign process_intf_32.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_continue;
    assign process_intf_32.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_start;
    assign process_intf_32.pin_stall = 1'b0;
    assign process_intf_32.pout_stall = 1'b0;
    assign process_intf_32.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_32;
    csv_file_dump pstatus_csv_dumper_32;
    df_process_monitor process_monitor_32;
    df_process_intf process_intf_33(clock,reset);
    assign process_intf_33.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_start;
    assign process_intf_33.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_ready;
    assign process_intf_33.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_done;
    assign process_intf_33.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_continue;
    assign process_intf_33.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_start;
    assign process_intf_33.pin_stall = 1'b0;
    assign process_intf_33.pout_stall = 1'b0;
    assign process_intf_33.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_33;
    csv_file_dump pstatus_csv_dumper_33;
    df_process_monitor process_monitor_33;
    df_process_intf process_intf_34(clock,reset);
    assign process_intf_34.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_start;
    assign process_intf_34.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_ready;
    assign process_intf_34.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_done;
    assign process_intf_34.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_continue;
    assign process_intf_34.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_start;
    assign process_intf_34.pin_stall = 1'b0;
    assign process_intf_34.pout_stall = 1'b0;
    assign process_intf_34.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_34;
    csv_file_dump pstatus_csv_dumper_34;
    df_process_monitor process_monitor_34;
    df_process_intf process_intf_35(clock,reset);
    assign process_intf_35.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.entry_proc_U0.ap_start;
    assign process_intf_35.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.entry_proc_U0.ap_ready;
    assign process_intf_35.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.entry_proc_U0.ap_done;
    assign process_intf_35.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.entry_proc_U0.ap_continue;
    assign process_intf_35.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.entry_proc_U0.ap_start;
    assign process_intf_35.pin_stall = 1'b0;
    assign process_intf_35.pout_stall = 1'b0;
    assign process_intf_35.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_35;
    csv_file_dump pstatus_csv_dumper_35;
    df_process_monitor process_monitor_35;
    df_process_intf process_intf_36(clock,reset);
    assign process_intf_36.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_start;
    assign process_intf_36.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_ready;
    assign process_intf_36.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_done;
    assign process_intf_36.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_continue;
    assign process_intf_36.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_start;
    assign process_intf_36.pin_stall = 1'b0;
    assign process_intf_36.pout_stall = 1'b0;
    assign process_intf_36.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_36;
    csv_file_dump pstatus_csv_dumper_36;
    df_process_monitor process_monitor_36;
    df_process_intf process_intf_37(clock,reset);
    assign process_intf_37.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_start;
    assign process_intf_37.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_ready;
    assign process_intf_37.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_done;
    assign process_intf_37.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_continue;
    assign process_intf_37.real_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_start;
    assign process_intf_37.pin_stall = 1'b0;
    assign process_intf_37.pout_stall = 1'b0;
    assign process_intf_37.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_37;
    csv_file_dump pstatus_csv_dumper_37;
    df_process_monitor process_monitor_37;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_fwd_fft.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_fwd_fft.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_fwd_fft.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_done;
    assign module_intf_6.ap_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_continue;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_done;
    assign module_intf_21.ap_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_continue;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_done;
    assign module_intf_22.ap_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_continue;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_done;
    assign module_intf_35.ap_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_continue;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;

    df_loop_intf df_loop_intf_1(clock,reset);
    assign df_loop_intf_1.body_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_start;
    assign df_loop_intf_1.body_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_ready;
    assign df_loop_intf_1.body_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_done;
    assign df_loop_intf_1.body_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.ap_continue;
    assign df_loop_intf_1.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_start;
    assign df_loop_intf_1.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_ready;
    assign df_loop_intf_1.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_done;
    assign df_loop_intf_1.loop_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.ap_continue;
    csv_file_dump df_loop_csv_dumper_1;
    df_loop_monitor df_loop_monitor_1;
    df_loop_intf df_loop_intf_2(clock,reset);
    assign df_loop_intf_2.body_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_start;
    assign df_loop_intf_2.body_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_ready;
    assign df_loop_intf_2.body_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_done;
    assign df_loop_intf_2.body_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_continue;
    assign df_loop_intf_2.loop_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_start;
    assign df_loop_intf_2.loop_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_ready;
    assign df_loop_intf_2.loop_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_done;
    assign df_loop_intf_2.loop_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.ap_continue;
    csv_file_dump df_loop_csv_dumper_2;
    df_loop_monitor df_loop_monitor_2;
    df_loop_intf df_loop_intf_3(clock,reset);
    assign df_loop_intf_3.body_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_start;
    assign df_loop_intf_3.body_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_ready;
    assign df_loop_intf_3.body_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_done;
    assign df_loop_intf_3.body_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_continue;
    assign df_loop_intf_3.loop_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_start;
    assign df_loop_intf_3.loop_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_ready;
    assign df_loop_intf_3.loop_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_done;
    assign df_loop_intf_3.loop_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.ap_continue;
    csv_file_dump df_loop_csv_dumper_3;
    df_loop_monitor df_loop_monitor_3;
    df_loop_intf df_loop_intf_4(clock,reset);
    assign df_loop_intf_4.body_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_start;
    assign df_loop_intf_4.body_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_ready;
    assign df_loop_intf_4.body_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_done;
    assign df_loop_intf_4.body_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ap_continue;
    assign df_loop_intf_4.loop_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_start;
    assign df_loop_intf_4.loop_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_ready;
    assign df_loop_intf_4.loop_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_done;
    assign df_loop_intf_4.loop_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.ap_continue;
    csv_file_dump df_loop_csv_dumper_4;
    df_loop_monitor df_loop_monitor_4;
    df_loop_intf df_loop_intf_5(clock,reset);
    assign df_loop_intf_5.body_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_start;
    assign df_loop_intf_5.body_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_ready;
    assign df_loop_intf_5.body_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_done;
    assign df_loop_intf_5.body_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.ap_continue;
    assign df_loop_intf_5.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_start;
    assign df_loop_intf_5.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_ready;
    assign df_loop_intf_5.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_done;
    assign df_loop_intf_5.loop_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.ap_continue;
    csv_file_dump df_loop_csv_dumper_5;
    df_loop_monitor df_loop_monitor_5;
    df_loop_intf df_loop_intf_6(clock,reset);
    assign df_loop_intf_6.body_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_start;
    assign df_loop_intf_6.body_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_ready;
    assign df_loop_intf_6.body_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_done;
    assign df_loop_intf_6.body_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_continue;
    assign df_loop_intf_6.loop_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_start;
    assign df_loop_intf_6.loop_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_ready;
    assign df_loop_intf_6.loop_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_done;
    assign df_loop_intf_6.loop_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.ap_continue;
    csv_file_dump df_loop_csv_dumper_6;
    df_loop_monitor df_loop_monitor_6;
    df_loop_intf df_loop_intf_7(clock,reset);
    assign df_loop_intf_7.body_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_start;
    assign df_loop_intf_7.body_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_ready;
    assign df_loop_intf_7.body_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_done;
    assign df_loop_intf_7.body_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_continue;
    assign df_loop_intf_7.loop_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_start;
    assign df_loop_intf_7.loop_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_ready;
    assign df_loop_intf_7.loop_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_done;
    assign df_loop_intf_7.loop_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.ap_continue;
    csv_file_dump df_loop_csv_dumper_7;
    df_loop_monitor df_loop_monitor_7;
    df_loop_intf df_loop_intf_8(clock,reset);
    assign df_loop_intf_8.body_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_start;
    assign df_loop_intf_8.body_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_ready;
    assign df_loop_intf_8.body_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_done;
    assign df_loop_intf_8.body_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ap_continue;
    assign df_loop_intf_8.loop_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_start;
    assign df_loop_intf_8.loop_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_ready;
    assign df_loop_intf_8.loop_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_done;
    assign df_loop_intf_8.loop_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.ap_continue;
    csv_file_dump df_loop_csv_dumper_8;
    df_loop_monitor df_loop_monitor_8;
    seq_loop_intf#(28) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state7;
    assign seq_loop_intf_1.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.pre_loop_state1 = 28'h0;
    assign seq_loop_intf_1.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state18;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state8;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state8;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state17;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(28) seq_loop_monitor_1;
    seq_loop_intf#(28) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state7;
    assign seq_loop_intf_2.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.pre_loop_state1 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state8;
    assign seq_loop_intf_2.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state28;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state18;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state18;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state27;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(28) seq_loop_monitor_2;
    seq_loop_intf#(28) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_3.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.pre_loop_state1 = 28'h0;
    assign seq_loop_intf_3.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.ap_ST_fsm_state28;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(28) seq_loop_monitor_3;
    seq_loop_intf#(11) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_4.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_4.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_fwd_fft.Row_Wise_Synch_U0.ap_ST_fsm_state11;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(11) seq_loop_monitor_4;
    seq_loop_intf#(14) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_5.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.pre_loop_state1 = 14'h0;
    assign seq_loop_intf_5.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_ST_fsm_state13;
    assign seq_loop_intf_5.post_states_valid = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.ap_ST_fsm_state12;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(14) seq_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_1.quit_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_1.loop_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_210_4_fu_260.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b0;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_2.quit_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_enable_reg_pp0_iter6;
    assign upc_loop_intf_2.loop_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_228_7_VITIS_LOOP_231_8_VITIS_LOOP_234_9_fu_270.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_3.quit_enable = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.loop_start = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_fwd_fft.Mem_Patch_Gen_U0.grp_Mem_Patch_Gen_Pipeline_VITIS_LOOP_220_6_fu_286.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b0;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_4.quit_enable = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.loop_start = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_fwd_fft.Col_Wise_Overlap_Gen_U0.grp_Col_Wise_Overlap_Gen_Pipeline_VITIS_LOOP_263_1_VITIS_LOOP_269_3_VITIS_LOOP_272_4_VITIS_LOOP_275_5_fu_116.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b0;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_done;
    assign upc_loop_intf_5.loop_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.stream_2_buf17_U0.ap_continue;
    assign upc_loop_intf_5.quit_at_end = 1'b0;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_VITIS_LOOP_40_1_fu_66.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_enable_reg_pp0_iter16;
    assign upc_loop_intf_7.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_enable_reg_pp0_iter16;
    assign upc_loop_intf_7.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_0_018_U0.grp_fft_stage_0_018_Pipeline_SKIP_X_fu_75.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_8.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_8.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_SKIP_X_fu_48.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_1_019_U0.grp_fft_stage_1_019_Pipeline_VITIS_LOOP_40_1_fu_61.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b0;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_10.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_10.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_2_020_U0.grp_fft_stage_2_020_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b0;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_12.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_12.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_3_021_U0.grp_fft_stage_3_021_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b0;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;
    upc_loop_intf#(1) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_14.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_14.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(1) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_4_022_U0.grp_fft_stage_4_022_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b0;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_enable_reg_pp0_iter17;
    assign upc_loop_intf_16.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_enable_reg_pp0_iter17;
    assign upc_loop_intf_16.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_SKIP_X_fu_46.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;
    upc_loop_intf#(1) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.fft_stage_5_023_U0.grp_fft_stage_5_023_Pipeline_VITIS_LOOP_40_1_fu_59.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b0;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(1) upc_loop_monitor_17;
    upc_loop_intf#(1) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.quit_state = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_18.quit_enable = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.loop_start = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_done;
    assign upc_loop_intf_18.loop_continue = AESL_inst_fwd_fft.FFT_R_U0.grp_dataflow_parent_loop_proc11_fu_112.dataflow_in_loop_VITIS_LOOP_91_1_U0.buf_2_stream24_U0.ap_continue;
    assign upc_loop_intf_18.quit_at_end = 1'b0;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(1) upc_loop_monitor_18;
    upc_loop_intf#(1) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.quit_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.quit_enable = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.loop_start = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_328_4_VITIS_LOOP_331_5_fu_152.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b0;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(1) upc_loop_monitor_19;
    upc_loop_intf#(1) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.quit_state = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.quit_block = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_start_enable = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.iter_end_enable = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_20.quit_enable = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.loop_start = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_fwd_fft.Row_Wise_Synch_U0.grp_Row_Wise_Synch_Pipeline_VITIS_LOOP_340_6_VITIS_LOOP_343_7_fu_161.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b0;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(1) upc_loop_monitor_20;
    upc_loop_intf#(1) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.quit_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.quit_enable = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.loop_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_done;
    assign upc_loop_intf_21.loop_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_gen_x_U0.ap_continue;
    assign upc_loop_intf_21.quit_at_end = 1'b0;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(1) upc_loop_monitor_21;
    upc_loop_intf#(1) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.quit_state = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_22.quit_enable = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_22.loop_start = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_done;
    assign upc_loop_intf_22.loop_continue = AESL_inst_fwd_fft.Transpose_U0.grp_dataflow_parent_loop_proc15_fu_82.dataflow_parent_loop_proc14_U0.dataflow_parent_loop_proc_U0.dataflow_in_loop_VITIS_LOOP_442_3_U0.ifmap_cons_y_U0.ap_continue;
    assign upc_loop_intf_22.quit_at_end = 1'b1;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(1) upc_loop_monitor_22;
    upc_loop_intf#(1) upc_loop_intf_23(clock,reset);
    assign upc_loop_intf_23.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_CS_fsm;
    assign upc_loop_intf_23.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_start;
    assign upc_loop_intf_23.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_ready;
    assign upc_loop_intf_23.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_done;
    assign upc_loop_intf_23.loop_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.stream_2_buf_U0.ap_continue;
    assign upc_loop_intf_23.quit_at_end = 1'b0;
    assign upc_loop_intf_23.finish = finish;
    csv_file_dump upc_loop_csv_dumper_23;
    upc_loop_monitor #(1) upc_loop_monitor_23;
    upc_loop_intf#(1) upc_loop_intf_24(clock,reset);
    assign upc_loop_intf_24.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_CS_fsm;
    assign upc_loop_intf_24.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_24.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_start;
    assign upc_loop_intf_24.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_ready;
    assign upc_loop_intf_24.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_VITIS_LOOP_40_1_fu_66.ap_done_int;
    assign upc_loop_intf_24.loop_continue = 1'b1;
    assign upc_loop_intf_24.quit_at_end = 1'b0;
    assign upc_loop_intf_24.finish = finish;
    csv_file_dump upc_loop_csv_dumper_24;
    upc_loop_monitor #(1) upc_loop_monitor_24;
    upc_loop_intf#(1) upc_loop_intf_25(clock,reset);
    assign upc_loop_intf_25.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_CS_fsm;
    assign upc_loop_intf_25.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_enable_reg_pp0_iter16;
    assign upc_loop_intf_25.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_enable_reg_pp0_iter16;
    assign upc_loop_intf_25.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_start;
    assign upc_loop_intf_25.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_ready;
    assign upc_loop_intf_25.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_0_0_U0.grp_fft_stage_0_0_Pipeline_SKIP_X_fu_75.ap_done_int;
    assign upc_loop_intf_25.loop_continue = 1'b1;
    assign upc_loop_intf_25.quit_at_end = 1'b1;
    assign upc_loop_intf_25.finish = finish;
    csv_file_dump upc_loop_csv_dumper_25;
    upc_loop_monitor #(1) upc_loop_monitor_25;
    upc_loop_intf#(1) upc_loop_intf_26(clock,reset);
    assign upc_loop_intf_26.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_CS_fsm;
    assign upc_loop_intf_26.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_26.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_26.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_26.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_start;
    assign upc_loop_intf_26.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_ready;
    assign upc_loop_intf_26.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_SKIP_X_fu_48.ap_done_int;
    assign upc_loop_intf_26.loop_continue = 1'b1;
    assign upc_loop_intf_26.quit_at_end = 1'b1;
    assign upc_loop_intf_26.finish = finish;
    csv_file_dump upc_loop_csv_dumper_26;
    upc_loop_monitor #(1) upc_loop_monitor_26;
    upc_loop_intf#(1) upc_loop_intf_27(clock,reset);
    assign upc_loop_intf_27.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_CS_fsm;
    assign upc_loop_intf_27.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_27.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_27.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_27.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_start;
    assign upc_loop_intf_27.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_ready;
    assign upc_loop_intf_27.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_1_0_U0.grp_fft_stage_1_0_Pipeline_VITIS_LOOP_40_1_fu_61.ap_done_int;
    assign upc_loop_intf_27.loop_continue = 1'b1;
    assign upc_loop_intf_27.quit_at_end = 1'b0;
    assign upc_loop_intf_27.finish = finish;
    csv_file_dump upc_loop_csv_dumper_27;
    upc_loop_monitor #(1) upc_loop_monitor_27;
    upc_loop_intf#(1) upc_loop_intf_28(clock,reset);
    assign upc_loop_intf_28.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_28.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_28.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_28.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_28.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_28.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_28.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_28.loop_continue = 1'b1;
    assign upc_loop_intf_28.quit_at_end = 1'b1;
    assign upc_loop_intf_28.finish = finish;
    csv_file_dump upc_loop_csv_dumper_28;
    upc_loop_monitor #(1) upc_loop_monitor_28;
    upc_loop_intf#(1) upc_loop_intf_29(clock,reset);
    assign upc_loop_intf_29.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_29.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_29.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_29.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_29.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_29.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_29.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_2_0_U0.grp_fft_stage_2_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_29.loop_continue = 1'b1;
    assign upc_loop_intf_29.quit_at_end = 1'b0;
    assign upc_loop_intf_29.finish = finish;
    csv_file_dump upc_loop_csv_dumper_29;
    upc_loop_monitor #(1) upc_loop_monitor_29;
    upc_loop_intf#(1) upc_loop_intf_30(clock,reset);
    assign upc_loop_intf_30.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_30.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_30.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_30.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_30.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_30.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_30.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_30.loop_continue = 1'b1;
    assign upc_loop_intf_30.quit_at_end = 1'b1;
    assign upc_loop_intf_30.finish = finish;
    csv_file_dump upc_loop_csv_dumper_30;
    upc_loop_monitor #(1) upc_loop_monitor_30;
    upc_loop_intf#(1) upc_loop_intf_31(clock,reset);
    assign upc_loop_intf_31.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_31.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_31.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_31.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_31.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_3_0_U0.grp_fft_stage_3_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_31.loop_continue = 1'b1;
    assign upc_loop_intf_31.quit_at_end = 1'b0;
    assign upc_loop_intf_31.finish = finish;
    csv_file_dump upc_loop_csv_dumper_31;
    upc_loop_monitor #(1) upc_loop_monitor_31;
    upc_loop_intf#(1) upc_loop_intf_32(clock,reset);
    assign upc_loop_intf_32.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_32.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_32.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_32.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_32.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_32.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_32.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_32.loop_continue = 1'b1;
    assign upc_loop_intf_32.quit_at_end = 1'b1;
    assign upc_loop_intf_32.finish = finish;
    csv_file_dump upc_loop_csv_dumper_32;
    upc_loop_monitor #(1) upc_loop_monitor_32;
    upc_loop_intf#(1) upc_loop_intf_33(clock,reset);
    assign upc_loop_intf_33.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_33.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_33.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_33.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_33.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_33.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_33.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_4_0_U0.grp_fft_stage_4_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_33.loop_continue = 1'b1;
    assign upc_loop_intf_33.quit_at_end = 1'b0;
    assign upc_loop_intf_33.finish = finish;
    csv_file_dump upc_loop_csv_dumper_33;
    upc_loop_monitor #(1) upc_loop_monitor_33;
    upc_loop_intf#(1) upc_loop_intf_34(clock,reset);
    assign upc_loop_intf_34.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_CS_fsm;
    assign upc_loop_intf_34.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_34.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter17;
    assign upc_loop_intf_34.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_enable_reg_pp0_iter17;
    assign upc_loop_intf_34.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_start;
    assign upc_loop_intf_34.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_ready;
    assign upc_loop_intf_34.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_SKIP_X_fu_50.ap_done_int;
    assign upc_loop_intf_34.loop_continue = 1'b1;
    assign upc_loop_intf_34.quit_at_end = 1'b1;
    assign upc_loop_intf_34.finish = finish;
    csv_file_dump upc_loop_csv_dumper_34;
    upc_loop_monitor #(1) upc_loop_monitor_34;
    upc_loop_intf#(1) upc_loop_intf_35(clock,reset);
    assign upc_loop_intf_35.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_CS_fsm;
    assign upc_loop_intf_35.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_35.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_35.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_35.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_start;
    assign upc_loop_intf_35.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_ready;
    assign upc_loop_intf_35.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.fft_stage_5_0_U0.grp_fft_stage_5_0_Pipeline_VITIS_LOOP_40_1_fu_63.ap_done_int;
    assign upc_loop_intf_35.loop_continue = 1'b1;
    assign upc_loop_intf_35.quit_at_end = 1'b0;
    assign upc_loop_intf_35.finish = finish;
    csv_file_dump upc_loop_csv_dumper_35;
    upc_loop_monitor #(1) upc_loop_monitor_35;
    upc_loop_intf#(1) upc_loop_intf_36(clock,reset);
    assign upc_loop_intf_36.cur_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_CS_fsm;
    assign upc_loop_intf_36.iter_start_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.iter_end_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.quit_state = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.iter_start_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.iter_end_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.quit_block = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.iter_start_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_36.iter_end_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_36.quit_enable = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_36.loop_start = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_start;
    assign upc_loop_intf_36.loop_ready = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_ready;
    assign upc_loop_intf_36.loop_done = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_done;
    assign upc_loop_intf_36.loop_continue = AESL_inst_fwd_fft.FFT_C_U0.grp_dataflow_parent_loop_proc12_fu_106.dataflow_in_loop_VITIS_LOOP_139_1_U0.buf_2_stream_U0.ap_continue;
    assign upc_loop_intf_36.quit_at_end = 1'b0;
    assign upc_loop_intf_36.finish = finish;
    csv_file_dump upc_loop_csv_dumper_36;
    upc_loop_monitor #(1) upc_loop_monitor_36;
    upc_loop_intf#(1) upc_loop_intf_37(clock,reset);
    assign upc_loop_intf_37.cur_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_CS_fsm;
    assign upc_loop_intf_37.iter_start_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.iter_end_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.quit_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.iter_start_block = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.iter_end_block = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.quit_block = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.iter_start_enable = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_37.iter_end_enable = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_37.quit_enable = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_37.loop_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_start;
    assign upc_loop_intf_37.loop_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_ready;
    assign upc_loop_intf_37.loop_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_done;
    assign upc_loop_intf_37.loop_continue = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_gen_y_U0.ap_continue;
    assign upc_loop_intf_37.quit_at_end = 1'b0;
    assign upc_loop_intf_37.finish = finish;
    csv_file_dump upc_loop_csv_dumper_37;
    upc_loop_monitor #(1) upc_loop_monitor_37;
    upc_loop_intf#(1) upc_loop_intf_38(clock,reset);
    assign upc_loop_intf_38.cur_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_CS_fsm;
    assign upc_loop_intf_38.iter_start_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.iter_end_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.quit_state = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.iter_start_block = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.iter_end_block = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.quit_block = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.iter_start_enable = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_38.iter_end_enable = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_38.quit_enable = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_38.loop_start = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_start;
    assign upc_loop_intf_38.loop_ready = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_ready;
    assign upc_loop_intf_38.loop_done = AESL_inst_fwd_fft.Mem_patch_Wr_U0.grp_dataflow_parent_loop_proc16_fu_70.dataflow_parent_loop_proc13_U0.dataflow_parent_loop_proc10_U0.dataflow_in_loop_VITIS_LOOP_471_3_U0.ifmap_vec_write_U0.grp_ifmap_vec_write_Pipeline_VITIS_LOOP_419_2_fu_107.ap_done_int;
    assign upc_loop_intf_38.loop_continue = 1'b1;
    assign upc_loop_intf_38.quit_at_end = 1'b0;
    assign upc_loop_intf_38.finish = finish;
    csv_file_dump upc_loop_csv_dumper_38;
    upc_loop_monitor #(1) upc_loop_monitor_38;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);
    fifo_csv_dumper_35 = new("./depth35.csv");
    cstatus_csv_dumper_35 = new("./chan_status35.csv");
    fifo_monitor_35 = new(fifo_csv_dumper_35,fifo_intf_35,cstatus_csv_dumper_35);
    fifo_csv_dumper_36 = new("./depth36.csv");
    cstatus_csv_dumper_36 = new("./chan_status36.csv");
    fifo_monitor_36 = new(fifo_csv_dumper_36,fifo_intf_36,cstatus_csv_dumper_36);
    fifo_csv_dumper_37 = new("./depth37.csv");
    cstatus_csv_dumper_37 = new("./chan_status37.csv");
    fifo_monitor_37 = new(fifo_csv_dumper_37,fifo_intf_37,cstatus_csv_dumper_37);
    fifo_csv_dumper_38 = new("./depth38.csv");
    cstatus_csv_dumper_38 = new("./chan_status38.csv");
    fifo_monitor_38 = new(fifo_csv_dumper_38,fifo_intf_38,cstatus_csv_dumper_38);
    fifo_csv_dumper_39 = new("./depth39.csv");
    cstatus_csv_dumper_39 = new("./chan_status39.csv");
    fifo_monitor_39 = new(fifo_csv_dumper_39,fifo_intf_39,cstatus_csv_dumper_39);
    fifo_csv_dumper_40 = new("./depth40.csv");
    cstatus_csv_dumper_40 = new("./chan_status40.csv");
    fifo_monitor_40 = new(fifo_csv_dumper_40,fifo_intf_40,cstatus_csv_dumper_40);
    fifo_csv_dumper_41 = new("./depth41.csv");
    cstatus_csv_dumper_41 = new("./chan_status41.csv");
    fifo_monitor_41 = new(fifo_csv_dumper_41,fifo_intf_41,cstatus_csv_dumper_41);
    fifo_csv_dumper_42 = new("./depth42.csv");
    cstatus_csv_dumper_42 = new("./chan_status42.csv");
    fifo_monitor_42 = new(fifo_csv_dumper_42,fifo_intf_42,cstatus_csv_dumper_42);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);
    pstall_csv_dumper_6 = new("./stalling6.csv");
    pstatus_csv_dumper_6 = new("./status6.csv");
    process_monitor_6 = new(pstall_csv_dumper_6,process_intf_6,pstatus_csv_dumper_6);
    pstall_csv_dumper_7 = new("./stalling7.csv");
    pstatus_csv_dumper_7 = new("./status7.csv");
    process_monitor_7 = new(pstall_csv_dumper_7,process_intf_7,pstatus_csv_dumper_7);
    pstall_csv_dumper_8 = new("./stalling8.csv");
    pstatus_csv_dumper_8 = new("./status8.csv");
    process_monitor_8 = new(pstall_csv_dumper_8,process_intf_8,pstatus_csv_dumper_8);
    pstall_csv_dumper_9 = new("./stalling9.csv");
    pstatus_csv_dumper_9 = new("./status9.csv");
    process_monitor_9 = new(pstall_csv_dumper_9,process_intf_9,pstatus_csv_dumper_9);
    pstall_csv_dumper_10 = new("./stalling10.csv");
    pstatus_csv_dumper_10 = new("./status10.csv");
    process_monitor_10 = new(pstall_csv_dumper_10,process_intf_10,pstatus_csv_dumper_10);
    pstall_csv_dumper_11 = new("./stalling11.csv");
    pstatus_csv_dumper_11 = new("./status11.csv");
    process_monitor_11 = new(pstall_csv_dumper_11,process_intf_11,pstatus_csv_dumper_11);
    pstall_csv_dumper_12 = new("./stalling12.csv");
    pstatus_csv_dumper_12 = new("./status12.csv");
    process_monitor_12 = new(pstall_csv_dumper_12,process_intf_12,pstatus_csv_dumper_12);
    pstall_csv_dumper_13 = new("./stalling13.csv");
    pstatus_csv_dumper_13 = new("./status13.csv");
    process_monitor_13 = new(pstall_csv_dumper_13,process_intf_13,pstatus_csv_dumper_13);
    pstall_csv_dumper_14 = new("./stalling14.csv");
    pstatus_csv_dumper_14 = new("./status14.csv");
    process_monitor_14 = new(pstall_csv_dumper_14,process_intf_14,pstatus_csv_dumper_14);
    pstall_csv_dumper_15 = new("./stalling15.csv");
    pstatus_csv_dumper_15 = new("./status15.csv");
    process_monitor_15 = new(pstall_csv_dumper_15,process_intf_15,pstatus_csv_dumper_15);
    pstall_csv_dumper_16 = new("./stalling16.csv");
    pstatus_csv_dumper_16 = new("./status16.csv");
    process_monitor_16 = new(pstall_csv_dumper_16,process_intf_16,pstatus_csv_dumper_16);
    pstall_csv_dumper_17 = new("./stalling17.csv");
    pstatus_csv_dumper_17 = new("./status17.csv");
    process_monitor_17 = new(pstall_csv_dumper_17,process_intf_17,pstatus_csv_dumper_17);
    pstall_csv_dumper_18 = new("./stalling18.csv");
    pstatus_csv_dumper_18 = new("./status18.csv");
    process_monitor_18 = new(pstall_csv_dumper_18,process_intf_18,pstatus_csv_dumper_18);
    pstall_csv_dumper_19 = new("./stalling19.csv");
    pstatus_csv_dumper_19 = new("./status19.csv");
    process_monitor_19 = new(pstall_csv_dumper_19,process_intf_19,pstatus_csv_dumper_19);
    pstall_csv_dumper_20 = new("./stalling20.csv");
    pstatus_csv_dumper_20 = new("./status20.csv");
    process_monitor_20 = new(pstall_csv_dumper_20,process_intf_20,pstatus_csv_dumper_20);
    pstall_csv_dumper_21 = new("./stalling21.csv");
    pstatus_csv_dumper_21 = new("./status21.csv");
    process_monitor_21 = new(pstall_csv_dumper_21,process_intf_21,pstatus_csv_dumper_21);
    pstall_csv_dumper_22 = new("./stalling22.csv");
    pstatus_csv_dumper_22 = new("./status22.csv");
    process_monitor_22 = new(pstall_csv_dumper_22,process_intf_22,pstatus_csv_dumper_22);
    pstall_csv_dumper_23 = new("./stalling23.csv");
    pstatus_csv_dumper_23 = new("./status23.csv");
    process_monitor_23 = new(pstall_csv_dumper_23,process_intf_23,pstatus_csv_dumper_23);
    pstall_csv_dumper_24 = new("./stalling24.csv");
    pstatus_csv_dumper_24 = new("./status24.csv");
    process_monitor_24 = new(pstall_csv_dumper_24,process_intf_24,pstatus_csv_dumper_24);
    pstall_csv_dumper_25 = new("./stalling25.csv");
    pstatus_csv_dumper_25 = new("./status25.csv");
    process_monitor_25 = new(pstall_csv_dumper_25,process_intf_25,pstatus_csv_dumper_25);
    pstall_csv_dumper_26 = new("./stalling26.csv");
    pstatus_csv_dumper_26 = new("./status26.csv");
    process_monitor_26 = new(pstall_csv_dumper_26,process_intf_26,pstatus_csv_dumper_26);
    pstall_csv_dumper_27 = new("./stalling27.csv");
    pstatus_csv_dumper_27 = new("./status27.csv");
    process_monitor_27 = new(pstall_csv_dumper_27,process_intf_27,pstatus_csv_dumper_27);
    pstall_csv_dumper_28 = new("./stalling28.csv");
    pstatus_csv_dumper_28 = new("./status28.csv");
    process_monitor_28 = new(pstall_csv_dumper_28,process_intf_28,pstatus_csv_dumper_28);
    pstall_csv_dumper_29 = new("./stalling29.csv");
    pstatus_csv_dumper_29 = new("./status29.csv");
    process_monitor_29 = new(pstall_csv_dumper_29,process_intf_29,pstatus_csv_dumper_29);
    pstall_csv_dumper_30 = new("./stalling30.csv");
    pstatus_csv_dumper_30 = new("./status30.csv");
    process_monitor_30 = new(pstall_csv_dumper_30,process_intf_30,pstatus_csv_dumper_30);
    pstall_csv_dumper_31 = new("./stalling31.csv");
    pstatus_csv_dumper_31 = new("./status31.csv");
    process_monitor_31 = new(pstall_csv_dumper_31,process_intf_31,pstatus_csv_dumper_31);
    pstall_csv_dumper_32 = new("./stalling32.csv");
    pstatus_csv_dumper_32 = new("./status32.csv");
    process_monitor_32 = new(pstall_csv_dumper_32,process_intf_32,pstatus_csv_dumper_32);
    pstall_csv_dumper_33 = new("./stalling33.csv");
    pstatus_csv_dumper_33 = new("./status33.csv");
    process_monitor_33 = new(pstall_csv_dumper_33,process_intf_33,pstatus_csv_dumper_33);
    pstall_csv_dumper_34 = new("./stalling34.csv");
    pstatus_csv_dumper_34 = new("./status34.csv");
    process_monitor_34 = new(pstall_csv_dumper_34,process_intf_34,pstatus_csv_dumper_34);
    pstall_csv_dumper_35 = new("./stalling35.csv");
    pstatus_csv_dumper_35 = new("./status35.csv");
    process_monitor_35 = new(pstall_csv_dumper_35,process_intf_35,pstatus_csv_dumper_35);
    pstall_csv_dumper_36 = new("./stalling36.csv");
    pstatus_csv_dumper_36 = new("./status36.csv");
    process_monitor_36 = new(pstall_csv_dumper_36,process_intf_36,pstatus_csv_dumper_36);
    pstall_csv_dumper_37 = new("./stalling37.csv");
    pstatus_csv_dumper_37 = new("./status37.csv");
    process_monitor_37 = new(pstall_csv_dumper_37,process_intf_37,pstatus_csv_dumper_37);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);

    df_loop_csv_dumper_1 = new("./df_loop_status1.csv");
    df_loop_monitor_1 = new(df_loop_intf_1,df_loop_csv_dumper_1);
    df_loop_csv_dumper_2 = new("./df_loop_status2.csv");
    df_loop_monitor_2 = new(df_loop_intf_2,df_loop_csv_dumper_2);
    df_loop_csv_dumper_3 = new("./df_loop_status3.csv");
    df_loop_monitor_3 = new(df_loop_intf_3,df_loop_csv_dumper_3);
    df_loop_csv_dumper_4 = new("./df_loop_status4.csv");
    df_loop_monitor_4 = new(df_loop_intf_4,df_loop_csv_dumper_4);
    df_loop_csv_dumper_5 = new("./df_loop_status5.csv");
    df_loop_monitor_5 = new(df_loop_intf_5,df_loop_csv_dumper_5);
    df_loop_csv_dumper_6 = new("./df_loop_status6.csv");
    df_loop_monitor_6 = new(df_loop_intf_6,df_loop_csv_dumper_6);
    df_loop_csv_dumper_7 = new("./df_loop_status7.csv");
    df_loop_monitor_7 = new(df_loop_intf_7,df_loop_csv_dumper_7);
    df_loop_csv_dumper_8 = new("./df_loop_status8.csv");
    df_loop_monitor_8 = new(df_loop_intf_8,df_loop_csv_dumper_8);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);
    upc_loop_csv_dumper_23 = new("./upc_loop_status23.csv");
    upc_loop_monitor_23 = new(upc_loop_intf_23,upc_loop_csv_dumper_23);
    upc_loop_csv_dumper_24 = new("./upc_loop_status24.csv");
    upc_loop_monitor_24 = new(upc_loop_intf_24,upc_loop_csv_dumper_24);
    upc_loop_csv_dumper_25 = new("./upc_loop_status25.csv");
    upc_loop_monitor_25 = new(upc_loop_intf_25,upc_loop_csv_dumper_25);
    upc_loop_csv_dumper_26 = new("./upc_loop_status26.csv");
    upc_loop_monitor_26 = new(upc_loop_intf_26,upc_loop_csv_dumper_26);
    upc_loop_csv_dumper_27 = new("./upc_loop_status27.csv");
    upc_loop_monitor_27 = new(upc_loop_intf_27,upc_loop_csv_dumper_27);
    upc_loop_csv_dumper_28 = new("./upc_loop_status28.csv");
    upc_loop_monitor_28 = new(upc_loop_intf_28,upc_loop_csv_dumper_28);
    upc_loop_csv_dumper_29 = new("./upc_loop_status29.csv");
    upc_loop_monitor_29 = new(upc_loop_intf_29,upc_loop_csv_dumper_29);
    upc_loop_csv_dumper_30 = new("./upc_loop_status30.csv");
    upc_loop_monitor_30 = new(upc_loop_intf_30,upc_loop_csv_dumper_30);
    upc_loop_csv_dumper_31 = new("./upc_loop_status31.csv");
    upc_loop_monitor_31 = new(upc_loop_intf_31,upc_loop_csv_dumper_31);
    upc_loop_csv_dumper_32 = new("./upc_loop_status32.csv");
    upc_loop_monitor_32 = new(upc_loop_intf_32,upc_loop_csv_dumper_32);
    upc_loop_csv_dumper_33 = new("./upc_loop_status33.csv");
    upc_loop_monitor_33 = new(upc_loop_intf_33,upc_loop_csv_dumper_33);
    upc_loop_csv_dumper_34 = new("./upc_loop_status34.csv");
    upc_loop_monitor_34 = new(upc_loop_intf_34,upc_loop_csv_dumper_34);
    upc_loop_csv_dumper_35 = new("./upc_loop_status35.csv");
    upc_loop_monitor_35 = new(upc_loop_intf_35,upc_loop_csv_dumper_35);
    upc_loop_csv_dumper_36 = new("./upc_loop_status36.csv");
    upc_loop_monitor_36 = new(upc_loop_intf_36,upc_loop_csv_dumper_36);
    upc_loop_csv_dumper_37 = new("./upc_loop_status37.csv");
    upc_loop_monitor_37 = new(upc_loop_intf_37,upc_loop_csv_dumper_37);
    upc_loop_csv_dumper_38 = new("./upc_loop_status38.csv");
    upc_loop_monitor_38 = new(upc_loop_intf_38,upc_loop_csv_dumper_38);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(fifo_monitor_35);
    sample_manager_inst.add_one_monitor(fifo_monitor_36);
    sample_manager_inst.add_one_monitor(fifo_monitor_37);
    sample_manager_inst.add_one_monitor(fifo_monitor_38);
    sample_manager_inst.add_one_monitor(fifo_monitor_39);
    sample_manager_inst.add_one_monitor(fifo_monitor_40);
    sample_manager_inst.add_one_monitor(fifo_monitor_41);
    sample_manager_inst.add_one_monitor(fifo_monitor_42);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(process_monitor_6);
    sample_manager_inst.add_one_monitor(process_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_8);
    sample_manager_inst.add_one_monitor(process_monitor_9);
    sample_manager_inst.add_one_monitor(process_monitor_10);
    sample_manager_inst.add_one_monitor(process_monitor_11);
    sample_manager_inst.add_one_monitor(process_monitor_12);
    sample_manager_inst.add_one_monitor(process_monitor_13);
    sample_manager_inst.add_one_monitor(process_monitor_14);
    sample_manager_inst.add_one_monitor(process_monitor_15);
    sample_manager_inst.add_one_monitor(process_monitor_16);
    sample_manager_inst.add_one_monitor(process_monitor_17);
    sample_manager_inst.add_one_monitor(process_monitor_18);
    sample_manager_inst.add_one_monitor(process_monitor_19);
    sample_manager_inst.add_one_monitor(process_monitor_20);
    sample_manager_inst.add_one_monitor(process_monitor_21);
    sample_manager_inst.add_one_monitor(process_monitor_22);
    sample_manager_inst.add_one_monitor(process_monitor_23);
    sample_manager_inst.add_one_monitor(process_monitor_24);
    sample_manager_inst.add_one_monitor(process_monitor_25);
    sample_manager_inst.add_one_monitor(process_monitor_26);
    sample_manager_inst.add_one_monitor(process_monitor_27);
    sample_manager_inst.add_one_monitor(process_monitor_28);
    sample_manager_inst.add_one_monitor(process_monitor_29);
    sample_manager_inst.add_one_monitor(process_monitor_30);
    sample_manager_inst.add_one_monitor(process_monitor_31);
    sample_manager_inst.add_one_monitor(process_monitor_32);
    sample_manager_inst.add_one_monitor(process_monitor_33);
    sample_manager_inst.add_one_monitor(process_monitor_34);
    sample_manager_inst.add_one_monitor(process_monitor_35);
    sample_manager_inst.add_one_monitor(process_monitor_36);
    sample_manager_inst.add_one_monitor(process_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(df_loop_monitor_1);
    sample_manager_inst.add_one_monitor(df_loop_monitor_2);
    sample_manager_inst.add_one_monitor(df_loop_monitor_3);
    sample_manager_inst.add_one_monitor(df_loop_monitor_4);
    sample_manager_inst.add_one_monitor(df_loop_monitor_5);
    sample_manager_inst.add_one_monitor(df_loop_monitor_6);
    sample_manager_inst.add_one_monitor(df_loop_monitor_7);
    sample_manager_inst.add_one_monitor(df_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_23);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_24);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_25);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_26);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_27);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_28);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_29);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_30);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_31);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_32);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_33);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_34);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_35);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_36);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_37);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_38);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
